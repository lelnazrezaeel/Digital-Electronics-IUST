** Profile: "SCHEMATIC1-2"  [ C:\USERS\SAEED\DESKTOP\pspicee\2-SCHEMATIC1-2.sim ] 

** Creating circuit file "2-SCHEMATIC1-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\2-SCHEMATIC1.net" 


.END
