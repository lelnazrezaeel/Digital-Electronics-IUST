** Profile: "SCHEMATIC1-3"  [ C:\USERS\SAEED\DESKTOP\pspicee\3-SCHEMATIC1-3.sim ] 

** Creating circuit file "3-SCHEMATIC1-3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\3-SCHEMATIC1.net" 


.END
